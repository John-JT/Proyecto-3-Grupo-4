`timescale 1ns / 1ps


module ALARMA_IMAGEN(
input bit_alarma,
input [9:0] Qh,
input [9:0] Qv,
input reloj,
input resetM,
output BIT_FUENTE5
    );
    
    
reg [255:0] data;
reg [8:0] addr_reg;
reg [7:0] SELEC_PX;
reg bit_fuente;

always@(*)begin
    SELEC_PX <= {Qh[7:0]};
    if (Qv[9:8] >= 3'd0 && Qv[9:8] < 3'd1)
    begin
        if (Qh[9:8] >= 3'd1 && Qh[9:8] < 3'd2)
            addr_reg <= {1'b0, Qv[7:0]};
        else    
            addr_reg <= 9'h1ff;
    end
    else
            addr_reg <= 9'h1ff;    
end

always@(posedge reloj)begin
        if (bit_alarma == 1'b1 && resetM == 1'b0)
        case (addr_reg)
        9'h000:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h001:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h002:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h003:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h004:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h005:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h006:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h007:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h008:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h009:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h00a:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h00b:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h00c:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h00d:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h00e:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h00f:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h010:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h011:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h012:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h013:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h014:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h015:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h016:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h017:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h018:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h019:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h01a:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h01b:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h01c:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h01d:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h01e:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h01f:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h020:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h021:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h022:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h023:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h024:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h025:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h026:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h027:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h028:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h029:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h02a:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h02b:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h02c:data <= 256'hfffffffffffffffffffffffffffffffffffffffffffffff8003fffcfffffffff;
        9'h02d:data <= 256'hfffffffff00000000000000100000000000001ffffffff000003ffc7ffffffff;
        9'h02e:data <= 256'hfffffffff00000000000000000000000000000fffffff8000000ff87ffffffff;
        9'h02f:data <= 256'hfffffffff00000000000000000000000000000ffffffe00000001f87ffffffff;
        9'h030:data <= 256'hfffffffff000000000000001fc000000000000ffffffc001ff800607ffffffff;
        9'h031:data <= 256'hfffffffff000000000000000ff000000000000ffffff000ffff80007ffffffff;
        9'h032:data <= 256'hfffffffff001fff001fff000ff8007ffffff00fffffc003fffff0007ffffffff;
        9'h033:data <= 256'hfffffffff00ffff001fffe00ff8007ffffff80fffff800ffffff8007ffffffff;
        9'h034:data <= 256'hfffffffff03ffff001ffff80ffc007ffffffe0fffff003ffffffc007ffffffff;
        9'h035:data <= 256'hfffffffff07ffff001ffffc0ffc007ffffffe0ffffe007fffffff007ffffffff;
        9'h036:data <= 256'hfffffffff0fffff001ffffe0ffc007fffffff0ffffc00ffffffff807ffffffff;
        9'h037:data <= 256'hfffffffff0fffff001fffff0ffc007fffffff0ffff801ffffffffc07ffffffff;
        9'h038:data <= 256'hfffffffff1fffff001fffff0ffc007fffffff0ffff003ffffffffc07ffffffff;
        9'h039:data <= 256'hfffffffff1fffff001fffff0ffc007fffffff8fffe003ffffffffe07ffffffff;
        9'h03a:data <= 256'hfffffffff1fffff001fffff8ffc007fffffff8fffc007fffffffff07ffffffff;
        9'h03b:data <= 256'hfffffffff3fffff001fffff8ffc007fffffff8fffc00ffffffffff07ffffffff;
        9'h03c:data <= 256'hfffffffff3fffff001fffff8ffc007fffffffcfff800ffffffffff87ffffffff;
        9'h03d:data <= 256'hfffffffff3fffff001fffffcffc007fffffffdfff001ffffffffff87ffffffff;
        9'h03e:data <= 256'hfffffffff3fffff001fffffdffc007fffffffffff001ffffffffffc3ffffffff;
        9'h03f:data <= 256'hfffffffffffffff001ffffffffc007ffffffffffe003ffffffffffc3ffffffff;
        9'h040:data <= 256'hfffffffffffffff001ffffffffc007ffffffffffe003ffffffffffe3ffffffff;
        9'h041:data <= 256'hfffffffffffffff001ffffffffc007ffffffffffc003ffffffffffe3ffffffff;
        9'h042:data <= 256'hfffffffffffffff001ffffffffc007ffffffffffc007fffffffffff3ffffffff;
        9'h043:data <= 256'hfffffffffffffff001ffffffffc007ffffff7fff8007fffffffffff3ffffffff;
        9'h044:data <= 256'hfffffffffffffff001ffffffffc007fffffe3fff8007fffffffffffbffffffff;
        9'h045:data <= 256'hfffffffffffffff001ffffffffc007fffffe3fff8007ffffffffffffffffffff;
        9'h046:data <= 256'hfffffffffffffff001ffffffffc007fffffe3fff000fffffffffffffffffffff;
        9'h047:data <= 256'hfffffffffffffff001ffffffffc007fffffe3fff000fffffffffffffffffffff;
        9'h048:data <= 256'hfffffffffffffff001ffffffffc007fffffc3fff000fffffffffffffffffffff;
        9'h049:data <= 256'hfffffffffffffff001ffffffffc007fffffc3fff000fffffffffffffffffffff;
        9'h04a:data <= 256'hfffffffffffffff001ffffffffc007fffffc3fff000fffffffffffffffffffff;
        9'h04b:data <= 256'hfffffffffffffff001ffffffffc007fffff83ffe000fffffffffffffffffffff;
        9'h04c:data <= 256'hfffffffffffffff001ffffffffc007ffffe03ffe001fffffffffffffffffffff;
        9'h04d:data <= 256'hfffffffffffffff001ffffffffc007ffff003ffe001fffffffffffffffffffff;
        9'h04e:data <= 256'hfffffffffffffff001ffffffffc0000000003ffe001fffffffffffffffffffff;
        9'h04f:data <= 256'hfffffffffffffff001ffffffffc0000000003ffe001fffffffffffffffffffff;
        9'h050:data <= 256'hfffffffffffffff001ffffffffc0000000003ffe001fffffffffffffffffffff;
        9'h051:data <= 256'hfffffffffffffff001ffffffffc0000000003ffe001fffffffffffffffffffff;
        9'h052:data <= 256'hfffffffffffffff001ffffffffc007ffff803ffe001fffffffffffffffffffff;
        9'h053:data <= 256'hfffffffffffffff001ffffffffc007fffff03ffe001fffffffffffffffffffff;
        9'h054:data <= 256'hfffffffffffffff001ffffffffc007fffff83ffe001fffffffffffffffffffff;
        9'h055:data <= 256'hfffffffffffffff001ffffffffc007fffffc3ffe001fffffffffffffffffffff;
        9'h056:data <= 256'hfffffffffffffff001ffffffffc007fffffc3ffe001fffffffffffffffffffff;
        9'h057:data <= 256'hfffffffffffffff001ffffffffc007fffffc3ffe001fffffffffffffffffffff;
        9'h058:data <= 256'hfffffffffffffff001ffffffffc007fffffc3ffe001fffffffffffffffffffff;
        9'h059:data <= 256'hfffffffffffffff001ffffffffc007fffffe3ffe000fffffffffffffffffffff;
        9'h05a:data <= 256'hfffffffffffffff001ffffffffc007fffffe3fff000fffffffffffffffffffff;
        9'h05b:data <= 256'hfffffffffffffff001ffffffffc007fffffe3fff000fffffffffffffffffffff;
        9'h05c:data <= 256'hfffffffffffffff001ffffffffc007fffffe7fff000fffffffffffffffffffff;
        9'h05d:data <= 256'hfffffffffffffff001ffffffffc007ffffffffff000fffffffffffffffffffff;
        9'h05e:data <= 256'hfffffffffffffff001ffffffffc007ffffffffff0007ffffffffffffffffffff;
        9'h05f:data <= 256'hfffffffffffffff001ffffffffc007ffffffffff8007ffffffffffffffffffff;
        9'h060:data <= 256'hfffffffffffffff001ffffffffc007ffffffffff8007ffffffffffffffffffff;
        9'h061:data <= 256'hfffffffffffffff001ffffffffc007ffffffffff8003ffffffffffffffffffff;
        9'h062:data <= 256'hfffffffffffffff001ffffffffc007ffffffffffc003ffffffffffffffffffff;
        9'h063:data <= 256'hfffffffffffffff001ffffffffc007ffffffffe7c003ffffffffffffffffffff;
        9'h064:data <= 256'hfffffffffffffff001ffffffffc007ffffffffc7e001fffffffffff8ffffffff;
        9'h065:data <= 256'hfffffffffffffff001ffffffffc007ffffffffc7e001fffffffffff1ffffffff;
        9'h066:data <= 256'hfffffffffffffff001ffffffffc007ffffffff87f000ffffffffffe1ffffffff;
        9'h067:data <= 256'hfffffffffffffff001ffffffffc007ffffffff8ff000ffffffffffe3ffffffff;
        9'h068:data <= 256'hfffffffffffffff001ffffffffc007ffffffff0ff8007fffffffffc7ffffffff;
        9'h069:data <= 256'hfffffffffffffff001ffffffffc007fffffffe0ffc003fffffffff87ffffffff;
        9'h06a:data <= 256'hfffffffffffffff001ffffffffc007fffffffe1ffe001fffffffff0fffffffff;
        9'h06b:data <= 256'hfffffffffffffff001ffffffffc007fffffffc1ffe000ffffffffe1fffffffff;
        9'h06c:data <= 256'hfffffffffffffff001ffffffffc007fffffff81fff0007fffffffc3fffffffff;
        9'h06d:data <= 256'hfffffffffffffff001ffffffffc007fffffff03fff8003fffffff87fffffffff;
        9'h06e:data <= 256'hfffffffffffffff001ffffffffc007ffffffe03fffc000ffffffe0ffffffffff;
        9'h06f:data <= 256'hfffffffffffffff001ffffffff8007ffffff807fffe0003fffffc1ffffffffff;
        9'h070:data <= 256'hffffffffffffffe000ffffffff8003fffffe007ffff8000fffff03ffffffffff;
        9'h071:data <= 256'hffffffffffffffc0007fffffff0000000000007ffffc0001fff007ffffffffff;
        9'h072:data <= 256'hffffffffffffff80003ffffffc000000000000fffffe000000001fffffffffff;
        9'h073:data <= 256'hffffffffffffc00000007fff00000000000000ffffff800000003fffffffffff;
        9'h074:data <= 256'hffffffffffffc00000007fff00000000000000ffffffe0000000ffffffffffff;
        9'h075:data <= 256'hffffffffffffe3e03000ffff3109180000f021fffffffc000007ffffffffffff;
        9'h076:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffe0007fffffffffffff;
        9'h077:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h078:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h079:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h07a:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h07b:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h07c:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h07d:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h07e:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h07f:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h080:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h081:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h082:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h083:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h084:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h085:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h086:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h087:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h088:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h089:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h08a:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h08b:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h08c:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h08d:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h08e:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h08f:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h090:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h091:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h092:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h093:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h094:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h095:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h096:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h097:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h098:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h099:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h09a:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h09b:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h09c:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h09d:data <= 256'hfffffffffffffffffffffffffffffffffbffffffffffffffffffffffffffffff;
        9'h09e:data <= 256'hfffffe00007fffffffffffffffffffffe3fffe3ffffffffc7fffffffffffffff;
        9'h09f:data <= 256'hfffffe00007fffffffffffffffffffff83fffe3ffffffffc7fffffffffffffff;
        9'h0a0:data <= 256'hfffffe7e3e7fffffffffffffffffffffe3fffc7ffffffffcffffffffffffffff;
        9'h0a1:data <= 256'hfffffefe3f3fffffffffffffffffffffe3fffcffffffffffffffffffffffffff;
        9'h0a2:data <= 256'hfffffffe3fbfffffffffffffffffffffe3fffdffffffffffffffffffffffffff;
        9'h0a3:data <= 256'hfffffffe3ffffffffffffffffffffffff3fffbffffffffffffffffffffffffff;
        9'h0a4:data <= 256'hfffffffe3ffffffffffffffffffffffff3ffffffffffffffffffffffffffffff;
        9'h0a5:data <= 256'hfffffffe3fffffffffffffffffffffffe3ffffffffffffffffffffffffffffff;
        9'h0a6:data <= 256'hfffffffe3fffc1fffc1ffe383fff03fff3fff03fffc1fffc7ffc0fffc0ffffff;
        9'h0a7:data <= 256'hfffffffe3fff087ff087fc303ffe20fff3ffc01fff3c0ff07ff007ff087fffff;
        9'h0a8:data <= 256'hfffffffe3ffe3c3fe3c7fe261ffcf87ff3ff8f8ffe3e3ff87ff3c3fe3e3fffff;
        9'h0a9:data <= 256'hfffffffe3ffe7e3fe7c3fe1f1ff8fc7ff3ff9fc7fe3e3ffc7fe7e3fe7f1fffff;
        9'h0aa:data <= 256'hfffffffe3ffc7e1fcfe7ff1f1ff1fc3ff3ff1fc7fe3f3ffc7fc7e3fc7f1fffff;
        9'h0ab:data <= 256'hfffffffe3ffc001fcfffff3f1ff1fe3ff3ff1fc3fe3e3ffc7fc7fffc7f0fffff;
        9'h0ac:data <= 256'hfffffffe3ffcffffcfffff3f1ff1fe3ff3ff3fe3fe3f3ffc7fc7fffc7f8fffff;
        9'h0ad:data <= 256'hfffffffe3ffcffffcfffff3f1ff1fe3ff3fe3fe3fe3e3ffc7fc7fffc7f8fffff;
        9'h0ae:data <= 256'hfffffffe3ffc7fffcfffff3f1ff1fe3ff3fe1fe3ff3e7ffc7fc7fffc7f8fffff;
        9'h0af:data <= 256'hfffffffe3ffc7fffc7fbff3f1ff1fe3ff3ff1fe3ff8cfffc7fc7fffc7f8fffff;
        9'h0b0:data <= 256'hfffffffe3ffc3fbfc7fbff3f1ff0fe3fe3ff1fe3ffa3fffc7fc3fffc7f8fffff;
        9'h0b1:data <= 256'hfffffffe3ffc1fbfc3f3ff3f1ff8fe3fe3ff0fc7fe7ffffc7fe3fbfc3f9fffff;
        9'h0b2:data <= 256'hfffffffc3ffe0f3fe0e7fe3f1ff87c7fe3ff8fc7fe7ffffc7fe0e3fe3f1fffff;
        9'h0b3:data <= 256'hfffffffc3fff007fe00ffe1f1ffc7cffe1ff878ffe001ffc7ff007fe1e3fffff;
        9'h0b4:data <= 256'hffffffe007ff00fff00ff80c07fe01ff80ffc01fff000ff01ff80fff807fffff;
        9'h0b5:data <= 256'hffffffffffffe3fffc3fffffffff87fffffff0ffff7fcffffffe3fffc1ffffff;
        9'h0b6:data <= 256'hfffffffffffffffffffffffffffffffffffffffffeffefffffffffffffffffff;
        9'h0b7:data <= 256'hfffffffffffffffffffffffffffffffffffffffffcffefffffffffffffffffff;
        9'h0b8:data <= 256'hfffffffffffffffffffffffffffffffffffffffffcffdfffffffffffffffffff;
        9'h0b9:data <= 256'hfffffffffffffffffffffffffffffffffffffffffc081fffffffffffffffffff;
        9'h0ba:data <= 256'hfffffffffffffffffffffffffffffffffffffffffe007fffffffffffffffffff;
        9'h0bb:data <= 256'hffffffffffffffffffffffffffffffffffffffffff81ffffffffffffffffffff;
        9'h0bc:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0bd:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0be:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0bf:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0c0:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0c1:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0c2:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffdfffffffffffffffff;
        9'h0c3:data <= 256'hffffffffe01fbfffffffffffffffffffffffefffffffff0fffffffffffffffff;
        9'h0c4:data <= 256'hffffffff00033fffffffffffffffffffffffe00003fffe0fffffffffffffffff;
        9'h0c5:data <= 256'hfffffffc07c03ffffffffffffffffffffffffc0000fffe0fffffffffffffffff;
        9'h0c6:data <= 256'hfffffff83ff83ffffffffffffffffffffffffe0fe03fff0fffffffffffffffff;
        9'h0c7:data <= 256'hfffffff07ffc1fffffffffffff7ffffffffffe0ff01fffffffffffffffffffff;
        9'h0c8:data <= 256'hffffffe0fffe1fffffffffffff3ffffffffffe0ff81fffffffffffffffffffff;
        9'h0c9:data <= 256'hffffffc1ffff1fffffffffffff3ffffffffffe0ffc0fffffffffffffffffffff;
        9'h0ca:data <= 256'hffffff83ffff1ffffffffffffe3ffffffffffe0ffc0fffffffffffffffffffff;
        9'h0cb:data <= 256'hffffff83ffff9ffffffffffffc3ffffffffffe0ffc0fffffffffffffffffffff;
        9'h0cc:data <= 256'hffffff03ffff9ffffffffffff83ffffffffffe0ffc0fffffffffffffffffffff;
        9'h0cd:data <= 256'hffffff07ffffdffffffffffff03ffffffffffe0ffc0fffffffffffffffffffff;
        9'h0ce:data <= 256'hffffff07fffffff803ffe003e001f801fffffe0ffc0fff0fff007ff003ffffff;
        9'h0cf:data <= 256'hfffffe07fffffff0c0ffc383c001f0e0fffffe0ffc1ffc0ffe183fe181ffffff;
        9'h0d0:data <= 256'hfffffe07ffffffe3f07fc7e3f83fe1f07ffffe0ff81ff00ff87c1fc3e0ffffff;
        9'h0d1:data <= 256'hfffffe07ffffffc7f83f8ff3f83fc3f87ffffe0ff03ffe0ff8fe0f87f0ffffff;
        9'h0d2:data <= 256'hfffffe0fffffff87fc1f8ff3f83fc3f87ffffe0fc07ffe0ff1fe0f87f0ffffff;
        9'h0d3:data <= 256'hfffffe0fffffff8ffc1f8ff3f83fc3f87ffffe0001ffff0fe1fe0f87f0ffffff;
        9'h0d4:data <= 256'hfffffe0fffffff0ffe0f87fbf83fc3f87ffffe0007ffff0fe1ff1f87f07fffff;
        9'h0d5:data <= 256'hfffffe0fffffff0ffe0f83fff83ffff83ffffe0f07ffff0fe1fffffff0ffffff;
        9'h0d6:data <= 256'hfffffe07ffffff0ffe0f807ff83fffc03ffffe0f03ffff0fc3ffffffc0ffffff;
        9'h0d7:data <= 256'hfffffe07fffffe0fff0fc03ff83fff003ffffe0f81ffff0fc3fffffe10ffffff;
        9'h0d8:data <= 256'hfffffe07fffffe0fff0fe00ff83ffc383ffffe0fc1ffff0fc1fffff830ffffff;
        9'h0d9:data <= 256'hfffffe07fffffe0fff0ff003f83ff0f83ffffe0fc0ffff0fc1ffffe1f0ffffff;
        9'h0da:data <= 256'hffffff07fffffe0fff0ffc01f83fe1f83ffffe0fe07fff0fc1ffffc3f0ffffff;
        9'h0db:data <= 256'hffffff03fffffe0fff0fff01f83fc3f83ffffe0ff03fff0fc1ffff87f0ffffff;
        9'h0dc:data <= 256'hffffff03ffffdf07ff0fbfc0f83fc3f83ffffe0ff83fff0fe0ffef87f07fffff;
        9'h0dd:data <= 256'hffffff81ffff9f07ff0fbfe0f83f83f83ffffe0ff81fff0fe0ffef07f07fffff;
        9'h0de:data <= 256'hffffffc1ffff9f03fe1fbff0f83f83f87ffffe0ffc0fff0fe07fcf07f07fffff;
        9'h0df:data <= 256'hffffffc0ffff3f83fe1f9ff0f83f83f83ffffe0ffe07ff0ff03f8f07f07fffff;
        9'h0e0:data <= 256'hffffffe03ffc7f81fc3f8ff1fc3d81e037fffe0ffe07ff0ff00e1f03c06fffff;
        9'h0e1:data <= 256'hfffffff00ff0ffc0fc7f87e1fc01c08007fffe07ff01fe0ff8003f80000fffff;
        9'h0e2:data <= 256'hfffffffc0001ffe030ff83c3fc03c0080ffffc03ff807c07fc007f80101fffff;
        9'h0e3:data <= 256'hffffffff0007fff801ff8007fe07e03c1fffe0007fc01001fe00ffc0783fffff;
        9'h0e4:data <= 256'hfffffffff03ffffe0ffffc3fffffffffffffffffffffffffff87ffffffffffff;
        9'h0e5:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0e6:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0e7:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0e8:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0e9:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0ea:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0eb:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0ec:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0ed:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0ee:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0ef:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0f0:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0f1:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0f2:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0f3:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0f4:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0f5:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0f6:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0f7:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0f8:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0f9:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0fa:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0fb:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0fc:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0fd:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0fe:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        9'h0ff:data <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
         
        default: data <= 256'd0;
        endcase
            else 
                data <= 256'd0;
    end
    always@(SELEC_PX, data, resetM , bit_alarma)begin
      if (bit_alarma == 1'b1 && resetM == 1'b0)
         case (SELEC_PX)
         8'b00000000: bit_fuente <= data[255];
         8'b00000001: bit_fuente <= data[254];
         8'b00000010: bit_fuente <= data[253];
         8'b00000011: bit_fuente <= data[252];
         8'b00000100: bit_fuente <= data[251];
         8'b00000101: bit_fuente <= data[250];
         8'b00000110: bit_fuente <= data[249];
         8'b00000111: bit_fuente <= data[248];
         8'b00001000: bit_fuente <= data[247];
         8'b00001001: bit_fuente <= data[246];
         8'b00001010: bit_fuente <= data[245];
         8'b00001011: bit_fuente <= data[244];
         8'b00001100: bit_fuente <= data[243];
         8'b00001101: bit_fuente <= data[242];
         8'b00001110: bit_fuente <= data[241];
         8'b00001111: bit_fuente <= data[240];
         8'b00010000: bit_fuente <= data[239];
         8'b00010001: bit_fuente <= data[238];
         8'b00010010: bit_fuente <= data[237];
         8'b00010011: bit_fuente <= data[236];
         8'b00010100: bit_fuente <= data[235];
         8'b00010101: bit_fuente <= data[234];
         8'b00010110: bit_fuente <= data[233];
         8'b00010111: bit_fuente <= data[232];
         8'b00011000: bit_fuente <= data[231];
         8'b00011001: bit_fuente <= data[230];
         8'b00011010: bit_fuente <= data[229];
         8'b00011011: bit_fuente <= data[228];
         8'b00011100: bit_fuente <= data[227];
         8'b00011101: bit_fuente <= data[226];
         8'b00011110: bit_fuente <= data[225];
         8'b00011111: bit_fuente <= data[224];
         8'b00100000: bit_fuente <= data[223];
         8'b00100001: bit_fuente <= data[222];
         8'b00100010: bit_fuente <= data[221];
         8'b00100011: bit_fuente <= data[220];
         8'b00100100: bit_fuente <= data[219];
         8'b00100101: bit_fuente <= data[218];
         8'b00100110: bit_fuente <= data[217];
         8'b00100111: bit_fuente <= data[216];
         8'b00101000: bit_fuente <= data[215];
         8'b00101001: bit_fuente <= data[214];
         8'b00101010: bit_fuente <= data[213];
         8'b00101011: bit_fuente <= data[212];
         8'b00101100: bit_fuente <= data[211];
         8'b00101101: bit_fuente <= data[210];
         8'b00101110: bit_fuente <= data[209];
         8'b00101111: bit_fuente <= data[208];
         8'b00110000: bit_fuente <= data[207];
         8'b00110001: bit_fuente <= data[206];
         8'b00110010: bit_fuente <= data[205];
         8'b00110011: bit_fuente <= data[204];
         8'b00110100: bit_fuente <= data[203];
         8'b00110101: bit_fuente <= data[202];
         8'b00110110: bit_fuente <= data[201];
         8'b00110111: bit_fuente <= data[200];
         8'b00111000: bit_fuente <= data[199];
         8'b00111001: bit_fuente <= data[198];
         8'b00111010: bit_fuente <= data[197];
         8'b00111011: bit_fuente <= data[196];
         8'b00111100: bit_fuente <= data[195];
         8'b00111101: bit_fuente <= data[194];
         8'b00111110: bit_fuente <= data[193];
         8'b00111111: bit_fuente <= data[192];
         8'b01000000: bit_fuente <= data[191];
         8'b01000001: bit_fuente <= data[190];
         8'b01000010: bit_fuente <= data[189];
         8'b01000011: bit_fuente <= data[188];
         8'b01000100: bit_fuente <= data[187];
         8'b01000101: bit_fuente <= data[186];
         8'b01000110: bit_fuente <= data[185];
         8'b01000111: bit_fuente <= data[184];
         8'b01001000: bit_fuente <= data[183];
         8'b01001001: bit_fuente <= data[182];
         8'b01001010: bit_fuente <= data[181];
         8'b01001011: bit_fuente <= data[180];
         8'b01001100: bit_fuente <= data[179];
         8'b01001101: bit_fuente <= data[178];
         8'b01001110: bit_fuente <= data[177];
         8'b01001111: bit_fuente <= data[176];
         8'b01010000: bit_fuente <= data[175];
         8'b01010001: bit_fuente <= data[174];
         8'b01010010: bit_fuente <= data[173];
         8'b01010011: bit_fuente <= data[172];
         8'b01010100: bit_fuente <= data[171];
         8'b01010101: bit_fuente <= data[170];
         8'b01010110: bit_fuente <= data[169];
         8'b01010111: bit_fuente <= data[168];
         8'b01011000: bit_fuente <= data[167];
         8'b01011001: bit_fuente <= data[166];
         8'b01011010: bit_fuente <= data[165];
         8'b01011011: bit_fuente <= data[164];
         8'b01011100: bit_fuente <= data[163];
         8'b01011101: bit_fuente <= data[162];
         8'b01011110: bit_fuente <= data[161];
         8'b01011111: bit_fuente <= data[160];
         8'b01100000: bit_fuente <= data[159];
         8'b01100001: bit_fuente <= data[158];
         8'b01100010: bit_fuente <= data[157];
         8'b01100011: bit_fuente <= data[156];
         8'b01100100: bit_fuente <= data[155];
         8'b01100101: bit_fuente <= data[154];
         8'b01100110: bit_fuente <= data[153];
         8'b01100111: bit_fuente <= data[152];
         8'b01101000: bit_fuente <= data[151];
         8'b01101001: bit_fuente <= data[150];
         8'b01101010: bit_fuente <= data[149];
         8'b01101011: bit_fuente <= data[148];
         8'b01101100: bit_fuente <= data[147];
         8'b01101101: bit_fuente <= data[146];
         8'b01101110: bit_fuente <= data[145];
         8'b01101111: bit_fuente <= data[144];
         8'b01110000: bit_fuente <= data[143];
         8'b01110001: bit_fuente <= data[142];
         8'b01110010: bit_fuente <= data[141];
         8'b01110011: bit_fuente <= data[140];
         8'b01110100: bit_fuente <= data[139];
         8'b01110101: bit_fuente <= data[138];
         8'b01110110: bit_fuente <= data[137];
         8'b01110111: bit_fuente <= data[136];
         8'b01111000: bit_fuente <= data[135];
         8'b01111001: bit_fuente <= data[134];
         8'b01111010: bit_fuente <= data[133];
         8'b01111011: bit_fuente <= data[132];
         8'b01111100: bit_fuente <= data[131];
         8'b01111101: bit_fuente <= data[130];
         8'b01111110: bit_fuente <= data[129];
         8'b01111111: bit_fuente <= data[128];         
         8'b10000000: bit_fuente <= data[127];
         8'b10000001: bit_fuente <= data[126];
         8'b10000010: bit_fuente <= data[125];
         8'b10000011: bit_fuente <= data[124];
         8'b10000100: bit_fuente <= data[123];
         8'b10000101: bit_fuente <= data[122];
         8'b10000110: bit_fuente <= data[121];
         8'b10000111: bit_fuente <= data[120];
         8'b10001000: bit_fuente <= data[119];
         8'b10001001: bit_fuente <= data[118];
         8'b10001010: bit_fuente <= data[117];
         8'b10001011: bit_fuente <= data[116];
         8'b10001100: bit_fuente <= data[115];
         8'b10001101: bit_fuente <= data[114];
         8'b10001110: bit_fuente <= data[113];
         8'b10001111: bit_fuente <= data[112];
         8'b10010000: bit_fuente <= data[111];
         8'b10010001: bit_fuente <= data[110];
         8'b10010010: bit_fuente <= data[109];
         8'b10010011: bit_fuente <= data[108];
         8'b10010100: bit_fuente <= data[107];
         8'b10010101: bit_fuente <= data[106];
         8'b10010110: bit_fuente <= data[105];
         8'b10010111: bit_fuente <= data[104];
         8'b10011000: bit_fuente <= data[103];
         8'b10011001: bit_fuente <= data[102];
         8'b10011010: bit_fuente <= data[101];
         8'b10011011: bit_fuente <= data[100];
         8'b10011100: bit_fuente <= data[99];
         8'b10011101: bit_fuente <= data[98];
         8'b10011110: bit_fuente <= data[97];
         8'b10011111: bit_fuente <= data[96];
         8'b10100000: bit_fuente <= data[95];
         8'b10100001: bit_fuente <= data[94];
         8'b10100010: bit_fuente <= data[93];
         8'b10100011: bit_fuente <= data[92];
         8'b10100100: bit_fuente <= data[91];
         8'b10100101: bit_fuente <= data[90];
         8'b10100110: bit_fuente <= data[89];
         8'b10100111: bit_fuente <= data[88];
         8'b10101000: bit_fuente <= data[87];
         8'b10101001: bit_fuente <= data[86];
         8'b10101010: bit_fuente <= data[85];
         8'b10101011: bit_fuente <= data[84];
         8'b10101100: bit_fuente <= data[83];
         8'b10101101: bit_fuente <= data[82];
         8'b10101110: bit_fuente <= data[81];
         8'b10101111: bit_fuente <= data[80];
         8'b10110000: bit_fuente <= data[79];
         8'b10110001: bit_fuente <= data[78];
         8'b10110010: bit_fuente <= data[77];
         8'b10110011: bit_fuente <= data[76];
         8'b10110100: bit_fuente <= data[75];
         8'b10110101: bit_fuente <= data[74];
         8'b10110110: bit_fuente <= data[73];
         8'b10110111: bit_fuente <= data[72];
         8'b10111000: bit_fuente <= data[71];
         8'b10111001: bit_fuente <= data[70];
         8'b10111010: bit_fuente <= data[69];
         8'b10111011: bit_fuente <= data[68];
         8'b10111100: bit_fuente <= data[67];
         8'b10111101: bit_fuente <= data[66];
         8'b10111110: bit_fuente <= data[65];
         8'b10111111: bit_fuente <= data[64];
         8'b11000000: bit_fuente <= data[63];
         8'b11000001: bit_fuente <= data[62];
         8'b11000010: bit_fuente <= data[61];
         8'b11000011: bit_fuente <= data[60];
         8'b11000100: bit_fuente <= data[59];
         8'b11000101: bit_fuente <= data[58];
         8'b11000110: bit_fuente <= data[57];
         8'b11000111: bit_fuente <= data[56];
         8'b11001000: bit_fuente <= data[55];
         8'b11001001: bit_fuente <= data[54];
         8'b11001010: bit_fuente <= data[53];
         8'b11001011: bit_fuente <= data[52];
         8'b11001100: bit_fuente <= data[51];
         8'b11001101: bit_fuente <= data[50];
         8'b11001110: bit_fuente <= data[49];
         8'b11001111: bit_fuente <= data[48];
         8'b11010000: bit_fuente <= data[47];
         8'b11010001: bit_fuente <= data[46];
         8'b11010010: bit_fuente <= data[45];
         8'b11010011: bit_fuente <= data[44];
         8'b11010100: bit_fuente <= data[43];
         8'b11010101: bit_fuente <= data[42];
         8'b11010110: bit_fuente <= data[41];
         8'b11010111: bit_fuente <= data[40];
         8'b11011000: bit_fuente <= data[39];
         8'b11011001: bit_fuente <= data[38];
         8'b11011010: bit_fuente <= data[37];
         8'b11011011: bit_fuente <= data[36];
         8'b11011100: bit_fuente <= data[35];
         8'b11011101: bit_fuente <= data[34];
         8'b11011110: bit_fuente <= data[33];
         8'b11011111: bit_fuente <= data[32];
         8'b11100000: bit_fuente <= data[31];
         8'b11100001: bit_fuente <= data[30];
         8'b11100010: bit_fuente <= data[29];
         8'b11100011: bit_fuente <= data[28];
         8'b11100100: bit_fuente <= data[27];
         8'b11100101: bit_fuente <= data[26];
         8'b11100110: bit_fuente <= data[25];
         8'b11100111: bit_fuente <= data[24];
         8'b11101000: bit_fuente <= data[23];
         8'b11101001: bit_fuente <= data[22];
         8'b11101010: bit_fuente <= data[21];
         8'b11101011: bit_fuente <= data[20];
         8'b11101100: bit_fuente <= data[19];
         8'b11101101: bit_fuente <= data[18];
         8'b11101110: bit_fuente <= data[17];
         8'b11101111: bit_fuente <= data[16];
         8'b11110000: bit_fuente <= data[15];
         8'b11110001: bit_fuente <= data[14];
         8'b11110010: bit_fuente <= data[13];
         8'b11110011: bit_fuente <= data[12];
         8'b11110100: bit_fuente <= data[11];
         8'b11110101: bit_fuente <= data[10];
         8'b11110110: bit_fuente <= data[9];
         8'b11110111: bit_fuente <= data[8];
         8'b11111000: bit_fuente <= data[7];
         8'b11111001: bit_fuente <= data[6];
         8'b11111010: bit_fuente <= data[5];
         8'b11111011: bit_fuente <= data[4];
         8'b11111100: bit_fuente <= data[3];
         8'b11111101: bit_fuente <= data[2];
         8'b11111110: bit_fuente <= data[1];
         8'b11111111: bit_fuente <= data[0];
          default:   bit_fuente <= 1'b0;
         endcase
         else
            bit_fuente <= 1'b0;
    end
    
    assign BIT_FUENTE5 = bit_fuente;
    
    
    
    
endmodule

